`ifndef YUU_INT_DEFINES_SVH
`define YUU_INT_DEFINES_SVH

  `ifndef YUU_MAX_INT_IDX
  `define YUU_MAX_INT_IDX 31
  `endif

`endif