`ifndef YUU_INT_TYPE_SVH
`define YUU_INT_TYPE_SVH

  typedef enum bit {
    POSEDGE,
    NEGEDGE 
    } yuu_int_severity_e;

`endif